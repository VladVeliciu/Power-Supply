* Netlist D:\College\4. year\Power Supplies\Project\Buck.psimsch *

.include "C:\Altair\Altair PSIM 2022.3\SPICElib\PSIM_SPICE.sub"

.tran 1.0e-006 1.0e-003 0  uic


.include "C:\Altair\Altair PSIM 2022.3\SPICElib\Diodes Inc\diode\Schottky diode models (Diodes Inc).txt"


SM_MOS1 1 2 3 0 SMM_MOS1 off
SMD_MOS1 2 1 2 1 SMDM_MOS1
.model SMM_MOS1 SW( Ron=1E-05 Roff=10meg Vt=0.5 Vh=0 )
.model SMDM_MOS1 SW( Ron=1E-05 Roff=10meg Vt=0 Vh=0 )
D_D1 0 4 B540C 
VI_IDIODE 2 4 0

L_L1 2 5 4.4E-05 Rser= 0.0002 IC= 0
VI_IL 5 6 0

R_R1 6 7 0.01
C_C1 7 8 0.0005 IC= 0
VI_ICap 8 0 0

E_VL VL 0 2 5 1
E_VTr VTr 0 2 1 1
VI_ITr 9 1 0

BV_ON1 3 0 V= IF( (V(10)>0.1), 1, 0 )
R_RL 11 0 1.65
VI_IOUT 6 11 0

V_VSQ 10 0 PULSE( 0 33 0 1E-07 1E-07 1.24E-05 5E-05 )
V_VDC1 12 0 DC 15
V_VTRI2 9 12 PULSE( 0 0.77 0.002 0.005 0.005 0 0.01 )
.save i(VI_IDIODE)
.save V(4)
.save i(VI_IL)
.save i(VI_ICap)
.save V(VL)
.save V(VTr)
.save i(VI_ITr)
.save i(VI_IOUT)
.save V(11)

* Matching PSIM probes to SPICE probes *
* IDIODE 	i(VI_IDIODE) *
* VDIODE 	V(4) *
* IL 	i(VI_IL) *
* ICap 	i(VI_ICap) *
* VL 	V(VL) *
* VTr 	V(VTr) *
* ITr 	i(VI_ITr) *
* IOUT 	i(VI_IOUT) *
* V2 	V(11) *

.end
